package mac_int32;

	interface mac_int32_ifc();
	endinterface

	(*synthesize*)
	module mkMAC_int32(mac_int32_ifc);
	endmodule


endpackage
